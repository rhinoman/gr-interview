Smith | Steve | steve@nowhere.com | Blue | 1979-05-02
Seldon | Hari | hari@foundation.net | Gray | 1988-01-01
Landale | Alis | alis@palma.net | Red | 1987-12-20
Burton | Levar | levar@burton.com | Red | 1957-02-16